Simultation of NMOS Inverter:

**inverter
VDD 2 0 5V
VIN 1 0 0V
R 3 2 1000
Mn 3 1 0 0 nMOD w=40u l=100u
.dc VIN 0v 5v .25v
.model nMOD nMOS(Vto=1 kp=25v
.plot dc V(3)
.probe
.end 