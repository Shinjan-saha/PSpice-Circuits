* C:\Users\SHINJAN SAHA\Documents\PSpice program\RTL.sch

* Schematics Version 9.1 - Web Update 1
* Tue Sep 05 12:52:00 2023



** Analysis setup **
.tran 0ms 1ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "RTL.net"
.INC "RTL.als"


.probe


.END
