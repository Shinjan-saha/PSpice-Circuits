* C:\Users\SHINJAN SAHA\Documents\PSpice program\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Tue Sep 05 12:10:28 2023



** Analysis setup **
.tran 0ns 1ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
